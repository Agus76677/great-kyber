module zetas_rom(
    input  wire [8:0] addr,
    output reg  [15:0] data
) ;
always @(*) begin
    case (addr)
        9'd0: data = 16'd1;
        9'd1: data = 16'd1;
        9'd2: data = 16'd1729;
        9'd3: data = 16'd1;
        9'd4: data = 16'd749;
        9'd5: data = 16'd1729;
        9'd6: data = 16'd40;
        9'd7: data = 16'd1;
        9'd8: data = 16'd2699;
        9'd9: data = 16'd749;
        9'd10: data = 16'd848;
        9'd11: data = 16'd1729;
        9'd12: data = 16'd2642;
        9'd13: data = 16'd40;
        9'd14: data = 16'd1432;
        9'd15: data = 16'd1;
        9'd16: data = 16'd797;
        9'd17: data = 16'd2699;
        9'd18: data = 16'd569;
        9'd19: data = 16'd749;
        9'd20: data = 16'd1062;
        9'd21: data = 16'd848;
        9'd22: data = 16'd69;
        9'd23: data = 16'd1729;
        9'd24: data = 16'd3136;
        9'd25: data = 16'd2642;
        9'd26: data = 16'd1746;
        9'd27: data = 16'd40;
        9'd28: data = 16'd1919;
        9'd29: data = 16'd1432;
        9'd30: data = 16'd2786;
        9'd31: data = 16'd1;
        9'd32: data = 16'd2240;
        9'd33: data = 16'd797;
        9'd34: data = 16'd936;
        9'd35: data = 16'd2699;
        9'd36: data = 16'd296;
        9'd37: data = 16'd569;
        9'd38: data = 16'd2882;
        9'd39: data = 16'd749;
        9'd40: data = 16'd3273;
        9'd41: data = 16'd1062;
        9'd42: data = 16'd1974;
        9'd43: data = 16'd848;
        9'd44: data = 16'd1990;
        9'd45: data = 16'd69;
        9'd46: data = 16'd1426;
        9'd47: data = 16'd1729;
        9'd48: data = 16'd1333;
        9'd49: data = 16'd3136;
        9'd50: data = 16'd450;
        9'd51: data = 16'd2642;
        9'd52: data = 16'd2447;
        9'd53: data = 16'd1746;
        9'd54: data = 16'd2794;
        9'd55: data = 16'd40;
        9'd56: data = 16'd3046;
        9'd57: data = 16'd1919;
        9'd58: data = 16'd821;
        9'd59: data = 16'd1432;
        9'd60: data = 16'd1853;
        9'd61: data = 16'd2786;
        9'd62: data = 16'd2094;
        9'd63: data = 16'd1;
        9'd64: data = 16'd2865;
        9'd65: data = 16'd2240;
        9'd66: data = 16'd2617;
        9'd67: data = 16'd797;
        9'd68: data = 16'd3040;
        9'd69: data = 16'd936;
        9'd70: data = 16'd1795;
        9'd71: data = 16'd2699;
        9'd72: data = 16'd2697;
        9'd73: data = 16'd296;
        9'd74: data = 16'd2474;
        9'd75: data = 16'd569;
        9'd76: data = 16'd2304;
        9'd77: data = 16'd2882;
        9'd78: data = 16'd1010;
        9'd79: data = 16'd749;
        9'd80: data = 16'd2009;
        9'd81: data = 16'd3273;
        9'd82: data = 16'd2681;
        9'd83: data = 16'd1062;
        9'd84: data = 16'd3253;
        9'd85: data = 16'd1974;
        9'd86: data = 16'd2868;
        9'd87: data = 16'd848;
        9'd88: data = 16'd2679;
        9'd89: data = 16'd1990;
        9'd90: data = 16'd2102;
        9'd91: data = 16'd69;
        9'd92: data = 16'd1274;
        9'd93: data = 16'd1426;
        9'd94: data = 16'd807;
        9'd95: data = 16'd1729;
        9'd96: data = 16'd33;
        9'd97: data = 16'd1333;
        9'd98: data = 16'd682;
        9'd99: data = 16'd3136;
        9'd100: data = 16'd2998;
        9'd101: data = 16'd450;
        9'd102: data = 16'd927;
        9'd103: data = 16'd2642;
        9'd104: data = 16'd2513;
        9'd105: data = 16'd2447;
        9'd106: data = 16'd3110;
        9'd107: data = 16'd1746;
        9'd108: data = 16'd2132;
        9'd109: data = 16'd2794;
        9'd110: data = 16'd1894;
        9'd111: data = 16'd40;
        9'd112: data = 16'd1414;
        9'd113: data = 16'd3046;
        9'd114: data = 16'd1481;
        9'd115: data = 16'd1919;
        9'd116: data = 16'd1756;
        9'd117: data = 16'd821;
        9'd118: data = 16'd1891;
        9'd119: data = 16'd1432;
        9'd120: data = 16'd1352;
        9'd121: data = 16'd1853;
        9'd122: data = 16'd2419;
        9'd123: data = 16'd2786;
        9'd124: data = 16'd2277;
        9'd125: data = 16'd2094;
        9'd126: data = 16'd452;
        9'd127: data = 16'd1;
        9'd128: data = 16'd939;
        9'd129: data = 16'd2865;
        9'd130: data = 16'd403;
        9'd131: data = 16'd2240;
        9'd132: data = 16'd2761;
        9'd133: data = 16'd2617;
        9'd134: data = 16'd561;
        9'd135: data = 16'd797;
        9'd136: data = 16'd2687;
        9'd137: data = 16'd3040;
        9'd138: data = 16'd1607;
        9'd139: data = 16'd936;
        9'd140: data = 16'd48;
        9'd141: data = 16'd1795;
        9'd142: data = 16'd1031;
        9'd143: data = 16'd2699;
        9'd144: data = 16'd992;
        9'd145: data = 16'd2697;
        9'd146: data = 16'd2443;
        9'd147: data = 16'd296;
        9'd148: data = 16'd1637;
        9'd149: data = 16'd2474;
        9'd150: data = 16'd2773;
        9'd151: data = 16'd569;
        9'd152: data = 16'd1651;
        9'd153: data = 16'd2304;
        9'd154: data = 16'd2935;
        9'd155: data = 16'd2882;
        9'd156: data = 16'd3050;
        9'd157: data = 16'd1010;
        9'd158: data = 16'd2954;
        9'd159: data = 16'd749;
        9'd160: data = 16'd892;
        9'd161: data = 16'd2009;
        9'd162: data = 16'd2237;
        9'd163: data = 16'd3273;
        9'd164: data = 16'd680;
        9'd165: data = 16'd2681;
        9'd166: data = 16'd735;
        9'd167: data = 16'd1062;
        9'd168: data = 16'd1847;
        9'd169: data = 16'd3253;
        9'd170: data = 16'd1874;
        9'd171: data = 16'd1974;
        9'd172: data = 16'd2662;
        9'd173: data = 16'd2868;
        9'd174: data = 16'd3220;
        9'd175: data = 16'd848;
        9'd176: data = 16'd641;
        9'd177: data = 16'd2679;
        9'd178: data = 16'd2186;
        9'd179: data = 16'd1990;
        9'd180: data = 16'd1041;
        9'd181: data = 16'd2102;
        9'd182: data = 16'd3010;
        9'd183: data = 16'd69;
        9'd184: data = 16'd1540;
        9'd185: data = 16'd1274;
        9'd186: data = 16'd1175;
        9'd187: data = 16'd1426;
        9'd188: data = 16'd756;
        9'd189: data = 16'd807;
        9'd190: data = 16'd2090;
        9'd191: data = 16'd1729;
        9'd192: data = 16'd2308;
        9'd193: data = 16'd33;
        9'd194: data = 16'd1026;
        9'd195: data = 16'd1333;
        9'd196: data = 16'd3312;
        9'd197: data = 16'd682;
        9'd198: data = 16'd1230;
        9'd199: data = 16'd3136;
        9'd200: data = 16'd1868;
        9'd201: data = 16'd2998;
        9'd202: data = 16'd2117;
        9'd203: data = 16'd450;
        9'd204: data = 16'd3096;
        9'd205: data = 16'd927;
        9'd206: data = 16'd1584;
        9'd207: data = 16'd2642;
        9'd208: data = 16'd733;
        9'd209: data = 16'd2513;
        9'd210: data = 16'd2775;
        9'd211: data = 16'd2447;
        9'd212: data = 16'd723;
        9'd213: data = 16'd3110;
        9'd214: data = 16'd757;
        9'd215: data = 16'd1746;
        9'd216: data = 16'd1626;
        9'd217: data = 16'd2132;
        9'd218: data = 16'd1219;
        9'd219: data = 16'd2794;
        9'd220: data = 16'd314;
        9'd221: data = 16'd1894;
        9'd222: data = 16'd780;
        9'd223: data = 16'd40;
        9'd224: data = 16'd941;
        9'd225: data = 16'd1414;
        9'd226: data = 16'd2804;
        9'd227: data = 16'd3046;
        9'd228: data = 16'd583;
        9'd229: data = 16'd1481;
        9'd230: data = 16'd2466;
        9'd231: data = 16'd1919;
        9'd232: data = 16'd952;
        9'd233: data = 16'd1756;
        9'd234: data = 16'd1029;
        9'd235: data = 16'd821;
        9'd236: data = 16'd1920;
        9'd237: data = 16'd1891;
        9'd238: data = 16'd1292;
        9'd239: data = 16'd1432;
        9'd240: data = 16'd3061;
        9'd241: data = 16'd1352;
        9'd242: data = 16'd1179;
        9'd243: data = 16'd1853;
        9'd244: data = 16'd2229;
        9'd245: data = 16'd2419;
        9'd246: data = 16'd1063;
        9'd247: data = 16'd2786;
        9'd248: data = 16'd2789;
        9'd249: data = 16'd2277;
        9'd250: data = 16'd885;
        9'd251: data = 16'd2094;
        9'd252: data = 16'd2156;
        9'd253: data = 16'd452;
        9'd254: data = 16'd1645;
        default: data = 16'd1;
    endcase
end
endmodule

module zetas_inv_rom(
    input  wire [8:0] addr,
    output reg  [15:0] data
) ;
always @(*) begin
    case (addr)
        9'd0: data = 16'd1;
        9'd1: data = 16'd1684;
        9'd2: data = 16'd2877;
        9'd3: data = 16'd1173;
        9'd4: data = 16'd1235;
        9'd5: data = 16'd2444;
        9'd6: data = 16'd1052;
        9'd7: data = 16'd540;
        9'd8: data = 16'd543;
        9'd9: data = 16'd2266;
        9'd10: data = 16'd910;
        9'd11: data = 16'd1100;
        9'd12: data = 16'd1476;
        9'd13: data = 16'd2150;
        9'd14: data = 16'd1977;
        9'd15: data = 16'd268;
        9'd16: data = 16'd1897;
        9'd17: data = 16'd2037;
        9'd18: data = 16'd1438;
        9'd19: data = 16'd1409;
        9'd20: data = 16'd2508;
        9'd21: data = 16'd2300;
        9'd22: data = 16'd1573;
        9'd23: data = 16'd2377;
        9'd24: data = 16'd1410;
        9'd25: data = 16'd863;
        9'd26: data = 16'd1848;
        9'd27: data = 16'd2746;
        9'd28: data = 16'd283;
        9'd29: data = 16'd525;
        9'd30: data = 16'd1915;
        9'd31: data = 16'd2388;
        9'd32: data = 16'd3289;
        9'd33: data = 16'd2549;
        9'd34: data = 16'd1435;
        9'd35: data = 16'd3015;
        9'd36: data = 16'd535;
        9'd37: data = 16'd2110;
        9'd38: data = 16'd1197;
        9'd39: data = 16'd1703;
        9'd40: data = 16'd1583;
        9'd41: data = 16'd2572;
        9'd42: data = 16'd219;
        9'd43: data = 16'd2606;
        9'd44: data = 16'd882;
        9'd45: data = 16'd554;
        9'd46: data = 16'd816;
        9'd47: data = 16'd2596;
        9'd48: data = 16'd687;
        9'd49: data = 16'd1745;
        9'd50: data = 16'd2402;
        9'd51: data = 16'd233;
        9'd52: data = 16'd2879;
        9'd53: data = 16'd1212;
        9'd54: data = 16'd331;
        9'd55: data = 16'd1461;
        9'd56: data = 16'd193;
        9'd57: data = 16'd2099;
        9'd58: data = 16'd2647;
        9'd59: data = 16'd17;
        9'd60: data = 16'd1996;
        9'd61: data = 16'd2303;
        9'd62: data = 16'd3296;
        9'd63: data = 16'd1021;
        9'd64: data = 16'd1600;
        9'd65: data = 16'd1239;
        9'd66: data = 16'd2522;
        9'd67: data = 16'd2573;
        9'd68: data = 16'd1903;
        9'd69: data = 16'd2154;
        9'd70: data = 16'd2055;
        9'd71: data = 16'd1789;
        9'd72: data = 16'd3260;
        9'd73: data = 16'd319;
        9'd74: data = 16'd1227;
        9'd75: data = 16'd2288;
        9'd76: data = 16'd1339;
        9'd77: data = 16'd1143;
        9'd78: data = 16'd650;
        9'd79: data = 16'd2688;
        9'd80: data = 16'd2481;
        9'd81: data = 16'd109;
        9'd82: data = 16'd461;
        9'd83: data = 16'd667;
        9'd84: data = 16'd1355;
        9'd85: data = 16'd1455;
        9'd86: data = 16'd76;
        9'd87: data = 16'd1482;
        9'd88: data = 16'd2267;
        9'd89: data = 16'd2594;
        9'd90: data = 16'd648;
        9'd91: data = 16'd2649;
        9'd92: data = 16'd56;
        9'd93: data = 16'd1092;
        9'd94: data = 16'd1320;
        9'd95: data = 16'd2437;
        9'd96: data = 16'd2580;
        9'd97: data = 16'd375;
        9'd98: data = 16'd2319;
        9'd99: data = 16'd279;
        9'd100: data = 16'd447;
        9'd101: data = 16'd394;
        9'd102: data = 16'd1025;
        9'd103: data = 16'd1678;
        9'd104: data = 16'd2760;
        9'd105: data = 16'd556;
        9'd106: data = 16'd855;
        9'd107: data = 16'd1692;
        9'd108: data = 16'd3033;
        9'd109: data = 16'd886;
        9'd110: data = 16'd632;
        9'd111: data = 16'd2337;
        9'd112: data = 16'd630;
        9'd113: data = 16'd2298;
        9'd114: data = 16'd1534;
        9'd115: data = 16'd3281;
        9'd116: data = 16'd2393;
        9'd117: data = 16'd1722;
        9'd118: data = 16'd289;
        9'd119: data = 16'd642;
        9'd120: data = 16'd2532;
        9'd121: data = 16'd2768;
        9'd122: data = 16'd712;
        9'd123: data = 16'd568;
        9'd124: data = 16'd1089;
        9'd125: data = 16'd2926;
        9'd126: data = 16'd464;
        9'd127: data = 16'd2390;
        9'd128: data = 16'd1;
        9'd129: data = 16'd2877;
        9'd130: data = 16'd1235;
        9'd131: data = 16'd1052;
        9'd132: data = 16'd543;
        9'd133: data = 16'd910;
        9'd134: data = 16'd1476;
        9'd135: data = 16'd1977;
        9'd136: data = 16'd1897;
        9'd137: data = 16'd1438;
        9'd138: data = 16'd2508;
        9'd139: data = 16'd1573;
        9'd140: data = 16'd1410;
        9'd141: data = 16'd1848;
        9'd142: data = 16'd283;
        9'd143: data = 16'd1915;
        9'd144: data = 16'd3289;
        9'd145: data = 16'd1435;
        9'd146: data = 16'd535;
        9'd147: data = 16'd1197;
        9'd148: data = 16'd1583;
        9'd149: data = 16'd219;
        9'd150: data = 16'd882;
        9'd151: data = 16'd816;
        9'd152: data = 16'd687;
        9'd153: data = 16'd2402;
        9'd154: data = 16'd2879;
        9'd155: data = 16'd331;
        9'd156: data = 16'd193;
        9'd157: data = 16'd2647;
        9'd158: data = 16'd1996;
        9'd159: data = 16'd3296;
        9'd160: data = 16'd1600;
        9'd161: data = 16'd2522;
        9'd162: data = 16'd1903;
        9'd163: data = 16'd2055;
        9'd164: data = 16'd3260;
        9'd165: data = 16'd1227;
        9'd166: data = 16'd1339;
        9'd167: data = 16'd650;
        9'd168: data = 16'd2481;
        9'd169: data = 16'd461;
        9'd170: data = 16'd1355;
        9'd171: data = 16'd76;
        9'd172: data = 16'd2267;
        9'd173: data = 16'd648;
        9'd174: data = 16'd56;
        9'd175: data = 16'd1320;
        9'd176: data = 16'd2580;
        9'd177: data = 16'd2319;
        9'd178: data = 16'd447;
        9'd179: data = 16'd1025;
        9'd180: data = 16'd2760;
        9'd181: data = 16'd855;
        9'd182: data = 16'd3033;
        9'd183: data = 16'd632;
        9'd184: data = 16'd630;
        9'd185: data = 16'd1534;
        9'd186: data = 16'd2393;
        9'd187: data = 16'd289;
        9'd188: data = 16'd2532;
        9'd189: data = 16'd712;
        9'd190: data = 16'd1089;
        9'd191: data = 16'd464;
        9'd192: data = 16'd1;
        9'd193: data = 16'd1235;
        9'd194: data = 16'd543;
        9'd195: data = 16'd1476;
        9'd196: data = 16'd1897;
        9'd197: data = 16'd2508;
        9'd198: data = 16'd1410;
        9'd199: data = 16'd283;
        9'd200: data = 16'd3289;
        9'd201: data = 16'd535;
        9'd202: data = 16'd1583;
        9'd203: data = 16'd882;
        9'd204: data = 16'd687;
        9'd205: data = 16'd2879;
        9'd206: data = 16'd193;
        9'd207: data = 16'd1996;
        9'd208: data = 16'd1600;
        9'd209: data = 16'd1903;
        9'd210: data = 16'd3260;
        9'd211: data = 16'd1339;
        9'd212: data = 16'd2481;
        9'd213: data = 16'd1355;
        9'd214: data = 16'd2267;
        9'd215: data = 16'd56;
        9'd216: data = 16'd2580;
        9'd217: data = 16'd447;
        9'd218: data = 16'd2760;
        9'd219: data = 16'd3033;
        9'd220: data = 16'd630;
        9'd221: data = 16'd2393;
        9'd222: data = 16'd2532;
        9'd223: data = 16'd1089;
        9'd224: data = 16'd1;
        9'd225: data = 16'd543;
        9'd226: data = 16'd1897;
        9'd227: data = 16'd1410;
        9'd228: data = 16'd3289;
        9'd229: data = 16'd1583;
        9'd230: data = 16'd687;
        9'd231: data = 16'd193;
        9'd232: data = 16'd1600;
        9'd233: data = 16'd3260;
        9'd234: data = 16'd2481;
        9'd235: data = 16'd2267;
        9'd236: data = 16'd2580;
        9'd237: data = 16'd2760;
        9'd238: data = 16'd630;
        9'd239: data = 16'd2532;
        9'd240: data = 16'd1;
        9'd241: data = 16'd1897;
        9'd242: data = 16'd3289;
        9'd243: data = 16'd687;
        9'd244: data = 16'd1600;
        9'd245: data = 16'd2481;
        9'd246: data = 16'd2580;
        9'd247: data = 16'd630;
        9'd248: data = 16'd1;
        9'd249: data = 16'd3289;
        9'd250: data = 16'd1600;
        9'd251: data = 16'd2580;
        9'd252: data = 16'd1;
        9'd253: data = 16'd1600;
        9'd254: data = 16'd1;
        default: data = 16'd1;
    endcase
end
endmodule

