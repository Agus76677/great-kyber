// Kyber NTT parameter definitions
localparam integer KYBER_Q        = 3329;
localparam integer KYBER_N        = 256;
localparam integer BARRETT_V      = 20159;
localparam integer BARRETT_SHIFT  = 26;
localparam integer BARRETT_ROUND  = 1 << 25;
localparam integer KYBER_N_INV    = 3316;
